countEasy
6
countNormal
6
countHard
6
maxEasy
1
maxNormal
1
maxHard
1
