countEasy
5
countNormal
5
countHard
5
maxEasy
1
maxNormal
1
maxHard
1
