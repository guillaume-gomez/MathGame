countEasy
4
countNormal
4
countHard
4
maxEasy
3
maxNormal
2
maxHard
1
