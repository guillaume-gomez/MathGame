countEasy
5
countNormal
5
countHard
5
maxEasy
4
maxNormal
4
maxHard
1
