countEasy
4
countNormal
4
countHard
4
maxEasy
4
maxNormal
4
maxHard
1
