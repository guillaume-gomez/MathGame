countEasy
7
countNormal
7
countHard
7
maxEasy
2
maxNormal
2
maxHard
1
