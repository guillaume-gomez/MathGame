countEasy
7countNormal
7countHard
7maxEasy
2maxNormal
2maxHard
1