countEasy
9countNormal
9countHard
9maxEasy
2maxNormal
2maxHard
1