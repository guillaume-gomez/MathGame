countEasy
7
countNormal
7
countHard
7
maxEasy
7
maxNormal
6
maxHard
6
