countEasy
13
countNormal
13
countHard
13
maxEasy
5
maxNormal
11
maxHard
8
