countEasy
6
countNormal
6
countHard
6
maxEasy
6
maxNormal
2
maxHard
2
