maxEasy
1
maxNormal
5
maxHard
1
