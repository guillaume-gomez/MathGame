countEasy
3
countNormal
3
countHard
3
maxEasy
3
maxNormal
2
maxHard
2
