countEasy
7
countNormal
7
countHard
7
maxEasy
6
maxNormal
6
maxHard
6
