countEasy
13
countNormal
13
countHard
13
maxEasy
5
maxNormal
13
maxHard
8
