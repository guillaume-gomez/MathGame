countEasy
2
countNormal
2
countHard
2
maxEasy
2
maxNormal
2
maxHard
1
