countEasy
7
countNormal
7
countHard
7
maxEasy
7
maxNormal
2
maxHard
2
