countEasy
2
countNormal
2
countHard
2
maxEasy
1
maxNormal
1
maxHard
1
