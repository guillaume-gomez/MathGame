countEasy
8
countNormal
8
countHard
8
maxEasy
2
maxNormal
2
maxHard
1
