countEasy
5
countNormal
5
countHard
5
maxEasy
3
maxNormal
2
maxHard
1
