countEasy
10countNormal
10countHard
10maxEasy
2maxNormal
2maxHard
1